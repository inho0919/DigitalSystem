--TB_HB_HA.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_HB_HA IS
END TB_HB_HA;

ARCHITECTURE HB OF TB_HB_HA IS
	COMPONENT HB_HA
		PORT(
			A, B : IN  BIT;
			D, U : OUT BIT
		);
	END COMPONENT;

	SIGNAL A, B : BIT := '0';
	SIGNAL D, U : BIT := '0';

BEGIN
	B <= '0', '1' AFTER 100 PS, '0' AFTER 200 PS, '1' AFTER 300 PS;
	A <= '0', '1' AFTER 200 PS;
	U_HB_HA : HB_HA
		PORT MAP(
			A => A,
			B => B,
			D => D,
			U => U
		);
END HB;
