--TB_HB_OR2.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_HB_OR2 IS
END TB_HB_OR2;

ARCHITECTURE HB OF TB_HB_OR2 IS
	COMPONENT HB_OR2
		PORT(
			A, B, C : IN  BIT;
			X    : OUT BIT
		);
	END COMPONENT;
	SIGNAL A : BIT := '0';
	SIGNAL B : BIT := '0';
	SIGNAL C : BIT := '0';
	SIGNAL X : BIT := '0';
BEGIN
	A <= '0', '1' AFTER 400 PS, '0' AFTER 800 PS;
	B <= '0', '1' AFTER 200 PS, '0' AFTER 400 PS, '1' AFTER 600 PS, '0' AFTER 800 PS;
	C <= '0', '1' AFTER 100 PS, '0' AFTER 200 PS, '1' AFTER 300 PS, '0' AFTER 400 PS, '1' AFTER 500 PS, '0' AFTER 600 PS, '1' AFTER 700 PS, '0' AFTER 800 PS;
	
	U_HB_OR2 : HB_OR2
		PORT MAP(
			A => A,
			B => B,
			C => C,
			X => X
		);
END HB;
