--TB_HB_OR2.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_HB_OR2 IS
END TB_HB_OR2;

ARCHITECTURE HB OF TB_HB_OR2 IS
	COMPONENT HB_OR2
		PORT(
			A, B : IN  BIT;
			X    : OUT BIT
		);
	END COMPONENT;
	SIGNAL A : BIT := '0';
	SIGNAL B : BIT := '0';
	SIGNAL X : BIT := '0';
BEGIN
	A <= '0', '1' AFTER 100 NS, '0' AFTER 300 NS, '1' AFTER 400 NS, '0' AFTER 500 NS;
	B <= '0', '1' AFTER 100 NS, '0' AFTER 200 NS, '1' AFTER 400 NS;
	U_HB_OR2 : HB_OR2
		PORT MAP(
			A => A,
			B => B,
			X => X
		);
END HB;
