-- TIMEBOMB_answer.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TIMEBOMB_answer IS
PORT(
	START 	 : IN  STD_LOGIC_VECTOR(0 DOWNTO 0);
	RESETN : IN STD_LOGIC;
	CLK_P : IN STD_LOGIC;
	CLK       : IN  STD_LOGIC;
	a, b, c, d, e, f, g : OUT STD_LOGIC;
	COUNT_OUT : BUFFER STD_LOGIC_VECTOR(0 TO 15); -- LED OUTPUT
	SEG_COM : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
	PIEZO : OUT STD_LOGIC
);
END TIMEBOMB_answer;

ARCHITECTURE HB OF TIMEBOMB_answer IS

	SIGNAL DECODE : STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL REG : STD_LOGIC;
	SIGNAL CNT : INTEGER RANGE 0 TO 2047;     
	SIGNAL LIMIT : INTEGER RANGE 0 TO 2047; 
	SIGNAL CNT_8BIT : STD_LOGIC_VECTOR(0 TO 15);
	SIGNAL HOLD : STD_LOGIC_VECTOR(0 DOWNTO 0);
	
	CONSTANT CNT_DO : INTEGER RANGE 0 TO 2047 := 1910;   
	CONSTANT CNT_MI : INTEGER RANGE 0 TO 2047 := 1516;
	CONSTANT CNT_SOL : INTEGER RANGE 0 TO 2047 := 1275; 
	CONSTANT CNT_HDO : INTEGER RANGE 0 TO 2047 := 955; 

BEGIN

SEG_COM <= "1";

PROCESS(START, RESETN, CLK)
	BEGIN
		IF START = 1 THEN
			IF RESETN = '0' THEN
				CNT_8BIT <= (OTHERS => '0');
			ELSIF CLK'EVENT AND CLK = '1' THEN
				IF CNT_8BIT = "11111111" THEN
					CNT_8BIT <= (OTHERS => '0');
				ELSE
					CNT_8BIT <= CNT_8BIT + 1;
				END IF;
			END IF;
		END IF;		
END PROCESS;

PROCESS(CLK) 
BEGIN     
	IF CNT_8BIT = "00001100" THEN   
		LIMIT <= CNT_DO;        
	ELSIF CNT_8BIT = "00001101" THEN    
		LIMIT <= CNT_MI;
   ELSIF CNT_8BIT = "00001110" THEN   
		LIMIT <= CNT_SOL;  
	ELSIF CNT_8BIT = "00001111" THEN    
		LIMIT <= CNT_HDO;   	
	ELSE 
		LIMIT <= 0;
	END IF; 
END PROCESS; 

PROCESS(RESETN, CLK_P) 
BEGIN  
   IF RESETN = '0' THEN 
	    CNT <= 0;     
	    REG <= '0';   
   ELSIF CLK_P'EVENT AND CLK_P = '1' THEN  
		IF CNT >= LIMIT THEN           
			CNT <= 0;         
			REG <= NOT REG;     
	    ELSE           
			CNT <= CNT + 1;      
	    END IF;  
   END IF; 
END PROCESS; 

PROCESS(CLK)
	BEGIN
		IF CNT_8BIT = "00001111" THEN
			COUNT_OUT <= "0000000000000001";
		ELSIF CNT_8BIT = "00001110" THEN
			COUNT_OUT <= "0000000000000010";
		ELSIF CNT_8BIT = "00001101" THEN
			COUNT_OUT <= "0000000000000100";	
		ELSIF CNT_8BIT = "00001100" THEN
			COUNT_OUT <= "0000000000001000";
		ELSIF CNT_8BIT = "00001011" THEN
			COUNT_OUT <= "0000000000010000";	
		ELSIF CNT_8BIT = "00001010" THEN
			COUNT_OUT <= "0000000000100000";
		ELSIF CNT_8BIT = "00001001" THEN
			COUNT_OUT <= "0000000001000000";
		ELSIF CNT_8BIT = "00001000" THEN
			COUNT_OUT <= "0000000010000000";
		ELSIF CNT_8BIT = "00000111" THEN
			COUNT_OUT <= "0000000100000000";
		ELSIF CNT_8BIT = "00000110" THEN
			COUNT_OUT <= "0000001000000000";
		ELSIF CNT_8BIT = "00000101" THEN
			COUNT_OUT <= "0000010000000000";
		ELSIF CNT_8BIT = "00000100" THEN
			COUNT_OUT <= "0000100000000000";
		ELSIF CNT_8BIT = "00000011" THEN
			COUNT_OUT <= "0001000000000000";
		ELSIF CNT_8BIT = "00000010" THEN
			COUNT_OUT <= "0010000000000000";
		ELSIF CNT_8BIT = "00000001" THEN
			COUNT_OUT <= "0100000000000000";
		ELSIF CNT_8BIT = "00000000" THEN
			COUNT_OUT <= "1000000000000000";
		ELSIF CNT_8BIT = "00010000" THEN
			COUNT_OUT <= "1010101001010101";
		ELSIF CNT_8BIT = "00010001" THEN
			COUNT_OUT <= "0101010110101010";	
		ELSIF CNT_8BIT = "00010010" THEN
			COUNT_OUT <= "1010101001010101";
		ELSIF CNT_8BIT = "00010011" THEN
			COUNT_OUT <= "0101010110101010";
		ELSIF CNT_8BIT = "00010100" THEN
			COUNT_OUT <= "1010101001010101";
		ELSIF CNT_8BIT = "00010101" THEN
			COUNT_OUT <= "0101010110101010";
		ELSE
			COUNT_OUT <= "1111111111111111";
		END IF;	
END PROCESS;
	
	
PROCESS(CLK)
	BEGIN
		CASE COUNT_OUT IS
			WHEN "1010101001010101" => DECODE <= "0000001";
			WHEN "0101010110101010" => DECODE <= "0110111";
			WHEN "1111111111111111" => DECODE <= "1111110"; 
			WHEN "0000000000000001" => DECODE <= "0110000"; 
			WHEN "0000000000000010" => DECODE <= "1101101"; 
			WHEN "0000000000000100" => DECODE <= "1111001"; 
			WHEN "0000000000001000" => DECODE <= "0110011"; 
			WHEN "0000000000010000" => DECODE <= "1011011"; 
			WHEN "0000000000100000" => DECODE <= "1011111"; 
			WHEN "0000000001000000" => DECODE <= "1110000"; 
			WHEN "0000000010000000" => DECODE <= "1111111"; 
			WHEN "0000000100000000" => DECODE <= "1111011"; 
			WHEN "0000001000000000" => DECODE <= "1110111"; 
			WHEN "0000010000000000" => DECODE <= "0011111"; 
			WHEN "0000100000000000" => DECODE <= "1001110"; 
			WHEN "0001000000000000" => DECODE <= "0111101"; 
			WHEN "0010000000000000" => DECODE <= "1001111"; 
			WHEN "0100000000000000" => DECODE <= "1000111"; 
			WHEN "1000000000000000" => DECODE <= "1100111"; 
			WHEN OTHERS => NULL;
		END CASE;
END PROCESS;

		
a <= DECODE(6);
b <= DECODE(5);
c <= DECODE(4);
d <= DECODE(3);
e <= DECODE(2);
f <= DECODE(1);
g <= DECODE(0);

PIEZO <= REG;

END HB;