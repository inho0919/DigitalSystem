--CLOCK.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CLOCK IS
	PORT(
		RESETN    : IN  STD_LOGIC;      -- RESET
		CLK       : IN  STD_LOGIC;      -- CLOCK 1Hz
		COUNT_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0) -- LED OUTPUT
	);
END CLOCK;

ARCHITECTURE HB OF CLOCK IS
	SIGNAL CNT_2BIT : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN
	PROCESS(RESETN, CLK)
	BEGIN
		IF RESETN = '0' THEN
			CNT_2BIT <= (OTHERS => '0');
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF CNT_2BIT = "11" THEN
				CNT_2BIT <= (OTHERS => '0');
			ELSE
				CNT_2BIT <= CNT_2BIT + 1;
			END IF;
		END IF;
	END PROCESS;
	COUNT_OUT <= CNT_2BIT;
END HB;