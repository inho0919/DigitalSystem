-- HB_OR2.VHD

ENTITY HB_OR2 IS
	PORT(
		A, B : IN BIT;
		X : OUT BIT
	);
END HB_OR2;

ARCHITECTURE HB OF HB_OR2 IS

BEGIN
	X <= A OR B;
END HB;